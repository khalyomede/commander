module commander

pub struct Argument {
    pub:
        name string
        description string
}
