module commander

fn (argument_list ArgumentList) is_filled() bool {
    return false
}
