module commander

pub type CommandFlag = Flag | TerminatingFlag
