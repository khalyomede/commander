module commander

pub struct Flag {
    pub:
        name string
        short_name string
        description string
}
